`include "define.v"
module wb(
	input clk,
	input rst
);

	always @ (posedge clk) begin
	end

	always @ (posedge clk) begin
	end
endmodule
